module FSMTester
(
		CLOCK_50,						//	On Board 50 MHz
		// Your inputs and outputs here
        KEY,
        SW,
		// The ports below are for the VGA output.  Do not change.
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK_N,						//	VGA BLANK
		VGA_SYNC_N,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B   						//	VGA Blue[9:0]
	);

	input			CLOCK_50;				//	50 MHz
	input   [9:0]   SW;
	input   [3:0]   KEY;

	// Do not change the following outputs
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK_N;				//	VGA BLANK
	output			VGA_SYNC_N;				//	VGA SYNC
	output	[9:0]	VGA_R;   				//	VGA Red[9:0]
	output	[9:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[9:0]	VGA_B;   				//	VGA Blue[9:0]
	
	wire resetn;
	assign resetn = KEY[0];
	
	// Create the colour, x, y and writeEn wires that are inputs to the controller.
	wire [2:0] gridColor, ezColor, normalColor, hardColor, clearColor;
	reg [2:0] color;
	reg [7:0] x;
	reg [6:0] y;
	
	wire [7: 0] gridXOut, ezXOut, normalXOut, hardXOut, clearXOut;
	wire [6: 0] gridYOut, ezYOut, normalYOut, hardYOut, clearYOut;
	
	
	wire grid, ez, normal, hard, inGame, clear;

	// Create an Instance of a VGA controller - there can be only one!
	// Define the number of colours as well as the initial background
	// image file (.MIF) for the controller.
	vga_adapter VGA(
			.resetn(resetn),
			.clock(CLOCK_50),
			.colour(color),
			.x(x),
			.y(y),
			.plot(SW[9]),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK_N),
			.VGA_SYNC(VGA_SYNC_N),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "160x120";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
		defparam VGA.BACKGROUND_IMAGE = "black.mif";
			
	// Put your code here. Your code should produce signals x,y,colour and writeEn/plot
	// for the VGA controller, in addition to any other functionality your design may require.
	 
	gameStateFSM gsfsm0(
		.clk(CLOCK_50),
		.resetn(KEY[0]),
		.go(~KEY[3:1]),
		.gameOver(SW[5]),
		.drawGrid(grid),
		.drawEZ(ez),
		.drawNORMAL(normal),
		.drawHARD(hard),
		.inGame(inGame),
		.clear(clear)
	);
	
	gridDrawer g0(
		.clk(CLOCK_50),
		.enable(grid),
		.resetn(KEY[0]),
		.colorOut(gridColor),
		.xOut(gridXOut),
		.yOut(gridYOut)
	);
	 
	numberDrawer d0(
		.numbers(64'b0000_1111_1110_1101_1100_1011_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001),
		.clk(CLOCK_50),
		.enable(ez),
		.resetn(KEY[0]),
		.colorOut(ezColor),
		.xOut(ezXOut),
		.yOut(ezYOut)
	);
	
	numberDrawer d1(
		.numbers(64'b0000_0001_0010_0011_0100_0101_0110_0111_1000_1001_1010_1011_1100_1101_1110_1111),
		.clk(CLOCK_50),
		.enable(normal),
		.resetn(KEY[0]),
		.colorOut(normalColor),
		.xOut(normalXOut),
		.yOut(normalYOut)
	);
	
	numberDrawer d2(
		.numbers(64'b0000_0101_0010_1011_0100_0001_0110_0011_1000_1001_1010_0111_1100_1101_1110_1111),
		.clk(CLOCK_50),
		.enable(hard),
		.resetn(KEY[0]),
		.colorOut(hardColor),
		.xOut(hardXOut),
		.yOut(hardYOut)
	);
	
	clear c0(
		.clk(CLOCK_50),
		.enable(clear),
		.resetn(KEY[0]),
		.colorOut(clearColor),
		.xOut(clearXOut),
		.yOut(clearYOut)
	);
	
	always@(*)
   begin
		if (grid == 1'b1)
			begin
				x = gridXOut;
				y = gridYOut;
				color = gridColor;
			end
		else if (ez == 1'b1)
			begin
				x = ezXOut;
				y = ezYOut;
				color = ezColor;
			end
		else if (normal == 1'b1)
			begin
				x = normalXOut;
				y = normalYOut;
				color = normalColor;
			end
		else if (hard == 1'b1)
			begin
				x = hardXOut;
				y = hardYOut;
				color = hardColor;
			end
		else if (clear == 1'b1)
			begin
				x = clearXOut;
				y = clearYOut;
				color = clearColor;
			end
		else
			begin
				x = 8'd0;
				y = 7'd0;
				color = 3'b000;
			end
	end
	
endmodule